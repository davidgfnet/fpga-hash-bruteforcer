-----------------------------------------------------------------------------------------------
--
--   E N T E R P O I N T   L T D
--
-----------------------------------------------------------------------------------------------
--
-- AUTHOR   : R FITZER
-- DATED    : 11/05/2012
--
-- COMMENTS : Cairnsmore 1 Test Program
--
--
-----------------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY UNISIM;
USE UNISIM.VCOMPONENTS.ALL;
--
ENTITY TOPLEVEL IS
PORT (
	-- 25MHz CLOCK FROM OSCILLATOR
	CLOCK_25MHZ			      : IN STD_LOGIC;
	--  CLOCKS FROM CLOCK GENERATOR
	CLK50					: IN STD_LOGIC;
	CLK100				: IN STD_LOGIC;
	CLK150				: IN STD_LOGIC;
	CLK200				: IN STD_LOGIC;

	CLOCKS1_2			: OUT STD_LOGIC;
	CLOCKS2_2			: OUT STD_LOGIC;
	CLOCKS3_2			: OUT STD_LOGIC;
	CLOCKS4_2			: OUT STD_LOGIC;
	-- ARRAY CLOCKS
	CLOCKS1_1			: OUT STD_LOGIC;
	CLOCKS2_1			: OUT STD_LOGIC;
	CLOCKS3_1			: OUT STD_LOGIC;
	CLOCKS4_1			: OUT STD_LOGIC;
	-- DIP SWITCHES
	SWITCH1				: IN STD_LOGIC;
	SWITCH2				: IN STD_LOGIC;
	SWITCH3				: IN STD_LOGIC;
	SWITCH4				: IN STD_LOGIC;
	SWITCH5				: IN STD_LOGIC;
	SWITCH6				: IN STD_LOGIC;
	SWITCH7				: IN STD_LOGIC;
	SWITCH8				: IN STD_LOGIC;
	-- POWER SUPPLY ENABLES
	EN_1V2_1				: OUT STD_LOGIC;
	EN_1V2_2				: OUT STD_LOGIC;
	EN_1V2_3				: OUT STD_LOGIC;
	EN_1V2_4				: OUT STD_LOGIC;
	ARRAY_3V3_EN		: OUT STD_LOGIC;
	-- SERIAL TO ARRAY FPGA 1
	USB1_1				: OUT STD_LOGIC;		-- TXD TO 	ARRAY 1
	USB1_2				: IN STD_LOGIC;		-- RXD FROM ARRAY 1
	-- SERIAL TO ARRAY FPGA 3
	USB3_1				: OUT STD_LOGIC;		-- TXD TO 	ARRAY 3
	USB3_2				: IN STD_LOGIC;		-- RXD FROM ARRAY 3
	-- JTAG DEDICATED - @ PORT 0
	USBC_0				: IN STD_LOGIC;		-- FTDI_TCK
	USBC_1				: IN STD_LOGIC;		-- FTDI_TDI
	USBC_2				: OUT STD_LOGIC;		-- FTDI_TDO
	USBC_3				: IN STD_LOGIC;		-- FTDI_TMS
	-- SPI DEDICATED - @ PORT 1
	USBC_8				: IN STD_LOGIC;		-- FTDI_SK
	USBC_9				: IN STD_LOGIC;		-- FTDI_DO
	USBC_10				: OUT STD_LOGIC;		-- FTDI_DI
	USBC_11				: IN STD_LOGIC;		-- FTDI_CS
	-- ICARUS STYLE PAIR @ PORT 1
	USBC_16				: IN STD_LOGIC;		-- FTDI_TXD
	USBC_17				: OUT STD_LOGIC;		-- FTDI_RXD
	-- ICARUS STYLE PAIR @ PORT 2
	USBC_24				: IN STD_LOGIC;		-- FTDI_TXD
	USBC_25				: OUT STD_LOGIC;		-- FTDI_RXD
	-- CLOCK GENERATOR
	CLK_SCLK          : OUT   STD_LOGIC;
	CLK_SDAT          : INOUT STD_LOGIC;
	-- JTAG DRIVE TO FPGA ARRAY ONLY WHEN SWITCH8 = 0
	JTAG_TCK				:  INOUT    STD_LOGIC;
	JTAG_TDI				:  INOUT    STD_LOGIC;
	JTAG_TDO				:  INOUT    STD_LOGIC;
	JTAG_TMS				:  INOUT    STD_LOGIC;
   
	USB1_5		      :  OUT      STD_LOGIC;		-- 1KHZ CLOCK
	USB2_5				:  OUT      STD_LOGIC;		-- 1KHZ CLOCK
	USB3_5				:  OUT      STD_LOGIC;		-- 1KHZ CLOCK
	USB4_5				:  OUT      STD_LOGIC;		-- 1KHZ CLOCK
   
	USB1_6		      :  OUT      STD_LOGIC;		-- RESET_N
	USB2_6				:  OUT      STD_LOGIC;		-- RESET_N
	USB3_6				:  OUT      STD_LOGIC;		-- RESET_N
	USB4_6				:  OUT      STD_LOGIC;		-- RESET_N
   
	USB1_7		      :  OUT      STD_LOGIC;		-- FREQUENCY_IS_100MHZ
	USB2_7				:  OUT      STD_LOGIC;		-- FREQUENCY_IS_100MHZ
	USB3_7				:  OUT      STD_LOGIC;		-- FREQUENCY_IS_100MHZ
	USB4_7				:  OUT      STD_LOGIC;		-- FREQUENCY_IS_100MHZ

	USB2_8				:  OUT      STD_LOGIC;		-- FREQUENCY_IS_100MHZ

   
	-- UPLINK 
	UP1	      		:  IN       STD_LOGIC;
	UP2			  		:  IN       STD_LOGIC;  
	UP3		   		:  IN       STD_LOGIC;
	UP4		   		:  IN       STD_LOGIC;
	-- DOWN LINK
	DOWN1	      		:  OUT      STD_LOGIC;
	DOWN2			  		:  OUT      STD_LOGIC;  
	DOWN3		   		:  OUT      STD_LOGIC;  
	DOWN4					:  OUT      STD_LOGIC;
   
   FAN_RPM1          :  IN       STD_LOGIC;
   FAN_RPM2          :  IN       STD_LOGIC;
   FAN_RPM3          :  IN       STD_LOGIC;
   FAN_RPM4          :  IN       STD_LOGIC;
   
	-- STATUS LED
	LED					:  OUT      STD_LOGIC
);
END TOPLEVEL;
--
ARCHITECTURE RTL OF TOPLEVEL IS
--
 	COMPONENT TX
	PORT(
		CLOCK				: IN STD_LOGIC;
		RESET				: IN STD_LOGIC;
		TX_ENABLE		: IN STD_LOGIC;
		TX_CHAR			: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		SERIAL_OUT  	: OUT STD_LOGIC;
		TX_BUSY     	: OUT STD_LOGIC
		);
	END COMPONENT;                                                     
--
 	COMPONENT RX
	PORT(
		CLOCK       	: IN STD_LOGIC;
		RESET				: IN STD_LOGIC;
		SERIAL_IN   	: IN STD_LOGIC;
		RX_CHAR			: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		RX_VALID	   	: OUT STD_LOGIC
		);
	END COMPONENT;                                                     
--
 	COMPONENT PULSE
	PORT (
		CLOCK       	: IN STD_LOGIC;
		RESET				: IN STD_LOGIC;
		TRIGGER   		: IN STD_LOGIC;
		STRETCHED  		: OUT STD_LOGIC
	);
	END COMPONENT;   
--	
COMPONENT FLASHER
    PORT ( CLOCK 			: IN  STD_LOGIC;
           RESET_N 		: IN  STD_LOGIC;
           COUNT 			: IN  INTEGER RANGE 0 TO 250000000;
			  FLASHOUT		: OUT	STD_LOGIC
			  );
END COMPONENT;

COMPONENT CLOCKGEN_CONTROLLER
  PORT( 
		CLOCK          	:  IN 	STD_LOGIC;
      RST_N             :  IN 	STD_LOGIC;
      CLK_SCLK          :  OUT   STD_LOGIC;
      CLK_SDAT          :  INOUT STD_LOGIC;
		IDT_SCLK      				:  OUT   STD_LOGIC;
		IDT_SDAT_OUT  				:  OUT   STD_LOGIC;  
		IDT_SDAT_OE   				:  OUT   STD_LOGIC;  
		IDT_SDAT_IN					:  OUT 	STD_LOGIC;
		IDT_EN_200KHZ				: OUT STD_LOGIC
      );                           
END COMPONENT;
--
COMPONENT LOOPBACK_TEST
	PORT(CLOCK_50MHZ 	      : IN  STD_LOGIC ;        
			RESET_N           : IN  STD_LOGIC ;    
			IO_TEST_BUS_IN    : IN  STD_LOGIC_VECTOR(1 TO 4);          
			IO_TEST_BUS_OUT   : OUT STD_LOGIC_VECTOR(1 TO 4);
			LOOPBACK_PASS	   : OUT STD_LOGIC  -- '1' = PASS
			);
END COMPONENT;
--
CONSTANT	MESSAGE_LENGTH	: INTEGER := 24;	
CONSTANT LOWERCASE_R		: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"72";
CONSTANT UPPERCASE_R		: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"52";
CONSTANT LOWERCASE_A		: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"61";
CONSTANT UPPERCASE_A		: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"41";
CONSTANT LOWERCASE_G		: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"67";
CONSTANT UPPERCASE_G		: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"47";
--
TYPE MESSAGESTATES IS ( IDLE, 
                        GETCHAR,
                        WAIT_BUSY,
                        WAIT_NOT_BUSY,
                        REPEAT
                        );
--
TYPE RXSTATES IS ( IDLE,
						GETCHAR,
						CHECK_R,
						CHECK_A,
						CHECK_G
						);							
--
SIGNAL RESET                  :  STD_LOGIC;
SIGNAL FLASH				      :  STD_LOGIC;
SIGNAL RESET_N				      :  STD_LOGIC;
SIGNAL CLOCK_100MHZ		      :  STD_LOGIC;
SIGNAL GCLOCKA				      :  STD_LOGIC;
--SIGNAL GCLOCKB				      :  STD_LOGIC;
--SIGNAL GCLOCKO				      :  STD_LOGIC;
SIGNAL GCLOCK				      :  STD_LOGIC;
SIGNAL SPI_DI				      :  STD_LOGIC;
SIGNAL SPI_SK				      :  STD_LOGIC;
SIGNAL SPI_CS				      :  STD_LOGIC;
SIGNAL SPI_DO				      :  STD_LOGIC;
SIGNAL SWITCH_STATE		      :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL IEN_1V2_1			      :  STD_LOGIC;
SIGNAL IEN_1V2_2			      :  STD_LOGIC;
SIGNAL IEN_1V2_3			      :  STD_LOGIC;
SIGNAL IEN_1V2_4			      :  STD_LOGIC;
SIGNAL IARRAY_3V3_EN		      :  STD_LOGIC;
SIGNAL LOOPIN1				      :  STD_LOGIC;
SIGNAL LOOPIN2				      :  STD_LOGIC;
SIGNAL LOOPIN3				      :  STD_LOGIC;
SIGNAL LOOPIN4				      :  STD_LOGIC;
SIGNAL LOOPOUT1			      :  STD_LOGIC;
SIGNAL LOOPOUT2			      :  STD_LOGIC;
SIGNAL LOOPOUT3			      :  STD_LOGIC;
SIGNAL LOOPOUT4			      :  STD_LOGIC;
SIGNAL LOOPBACK_PASS		      :  STD_LOGIC;
SIGNAL CLOCK_STOP			      :  STD_LOGIC;
SIGNAL TOGGLE_1KHZ            :  STD_LOGIC;
SIGNAL CLOCK_1KHZ             :  STD_LOGIC;
SIGNAL CLOCK_DIVIDE_COUNTER   :  INTEGER RANGE 0 TO 25000;
SIGNAL FREQUENCY_IS_100MHZ    :  STD_LOGIC;
SIGNAL COUNTER_100MS          :  INTEGER RANGE 0 TO 24999999;
SIGNAL COUNTER_100MS_TICK     :  STD_LOGIC;
SIGNAL POWER_STARTUP_N        :  STD_LOGIC_VECTOR( 5 DOWNTO 0);
SIGNAL OP_CLK_PHASE           :  STD_LOGIC_VECTOR( 3 DOWNTO 0);
SIGNAL FREQUENCY_IS_50MHZ     :  STD_LOGIC;
SIGNAL RESET_COUNT            :  STD_LOGIC_VECTOR( 7 DOWNTO 0);
SIGNAL RESET_FROM_COUNT       :  STD_LOGIC;
SIGNAL FAN_COUNTER1           :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL FAN_COUNTER2           :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL FAN_COUNTER3           :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL FAN_COUNTER4           :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL FAN_COUNTER1_STORED    :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL FAN_COUNTER2_STORED    :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL FAN_COUNTER3_STORED    :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL FAN_COUNTER4_STORED    :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL TICK_1SEC              :  STD_LOGIC;
SIGNAL TICK_COUNTER           :  INTEGER RANGE 0 TO 24999999;
SIGNAL FAN_RPM1_SHIFT         :  STD_LOGIC_VECTOR( 3 DOWNTO 0);
SIGNAL FAN_RPM2_SHIFT         :  STD_LOGIC_VECTOR( 3 DOWNTO 0);
SIGNAL FAN_RPM3_SHIFT         :  STD_LOGIC_VECTOR( 3 DOWNTO 0);
SIGNAL FAN_RPM4_SHIFT         :  STD_LOGIC_VECTOR( 3 DOWNTO 0);
SIGNAL FAN1_IS_OK             :  STD_LOGIC;
SIGNAL FAN2_IS_OK             :  STD_LOGIC;
SIGNAL FAN3_IS_OK             :  STD_LOGIC;
SIGNAL FAN4_IS_OK             :  STD_LOGIC;
SIGNAL FAN_IS_RUNNING         :  STD_LOGIC;
--
BEGIN

MAKE_A_RESET : PROCESS(SWITCH1,CLOCK_25MHZ)
BEGIN
IF (SWITCH1 = '1') THEN
   RESET_COUNT          <= X"00";
   RESET_FROM_COUNT     <= '1';
   
ELSIF (CLOCK_25MHZ'EVENT  AND CLOCK_25MHZ='1') THEN
   IF (RESET_COUNT = X"34") THEN
      RESET_COUNT          <= X"34";   
      RESET_FROM_COUNT     <= '0';
   ELSE
      RESET_COUNT          <= RESET_COUNT + 1;
      RESET_FROM_COUNT     <= '1';
   END IF;  
    
END IF;
END PROCESS MAKE_A_RESET;


RST : PROCESS(SWITCH1,RESET_FROM_COUNT,CLK50)
BEGIN
IF (RESET_FROM_COUNT = '1') THEN
   RESET_N <= '0';
ELSIF (CLK50'EVENT  AND CLK50='1') THEN
   RESET_N <= '1';
END IF;
END PROCESS RST;

RESET <= NOT RESET_N;


--
-- CONFIDENCE TICKER
--
TCK : FLASHER
    PORT MAP ( 
		CLOCK 		=> GCLOCK,
      RESET_N 		=> RESET_N,
      COUNT 		=> 12500000,
		FLASHOUT		=> FLASH
		);
--
CGEN : CLOCKGEN_CONTROLLER
  PORT MAP( 
		CLOCK				=> CLOCK_25MHZ,
      RST_N       	=> RESET_N,
      CLK_SCLK    	=> CLK_SCLK,
      CLK_SDAT    	=> CLK_SDAT,
		IDT_SCLK     	=> OPEN,   
		IDT_SDAT_OUT 	=> OPEN,
		IDT_SDAT_OE  	=> OPEN, 
		IDT_SDAT_IN	 	=> OPEN,
		IDT_EN_200KHZ  => OPEN
      );   
--
-- FLASH SPARTAN3 LED
--
-- ROUTE 100MHZ CLOCK TO ARRAY FPGA'S

OPCLKS : PROCESS(POWER_STARTUP_N,GCLOCK)
BEGIN
IF (POWER_STARTUP_N(5) = '1') THEN
   OP_CLK_PHASE   <= "0101";
   
   CLOCKS1_1	   <= '0';
   CLOCKS2_1	   <= '0';
   CLOCKS3_1	   <= '0';
   CLOCKS4_1	   <= '0';
   CLOCKS1_2	   <= '1';
   CLOCKS2_2	   <= '1';
   USB2_8         <= '1';
   CLOCKS3_2	   <= '1';
   CLOCKS4_2	   <= '1';
   
ELSIF (GCLOCK'EVENT  AND GCLOCK='1') THEN

   OP_CLK_PHASE( 3 DOWNTO 0)  <= OP_CLK_PHASE(2 DOWNTO 0) & OP_CLK_PHASE(3);

   CLOCKS1_1	   <= OP_CLK_PHASE(0);
   CLOCKS2_1	   <= OP_CLK_PHASE(1);
   CLOCKS3_1	   <= OP_CLK_PHASE(2);
   CLOCKS4_1	   <= OP_CLK_PHASE(3);
   
	CLOCKS1_2		<= OP_CLK_PHASE(1);
	CLOCKS2_2		<= OP_CLK_PHASE(2);
   USB2_8         <= OP_CLK_PHASE(2);
	CLOCKS3_2		<= OP_CLK_PHASE(3);
	CLOCKS4_2		<= OP_CLK_PHASE(0);
   
   
   
END IF;
END PROCESS OPCLKS;




--
-- Stop the clocks when we program!!
-- S = 1 = Stopped
--
-- 6 5
-- 0 0 - 50
-- 0 1 - 100
-- 1 0 - 150
-- 1 1 - 200
--
   BGMUX_50_100 : BUFGMUX
   port map (
      O 	=>	GCLOCKA,    
      I0 =>	CLK100,
      I1 => CLK200,  
      S 	=> SWITCH5
   );
--
   BGMUX_ON_OFF : BUFGMUX
   port map (
      O 	=>	GCLOCK,    
      I0 =>	GCLOCKA,
      I1 => '0',  
      S 	=> CLOCK_STOP
   );
--
SPI_ACCESS_inst : SPI_ACCESS
   generic map (
      SIM_DELAY_TYPE => "SCALED",
      SIM_DEVICE => "3S50AN",
      SIM_FACTORY_ID => X"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
      SIM_MEM_FILE => "NONE",
      SIM_USER_ID => X"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
   port map (
      MISO 	=> SPI_DI,
      CLK 	=> SPI_SK,
      CSB 	=> SPI_CS,
      MOSI 	=> SPI_DO
   );
--
-- JTAG Signals driven from USB Port 0 when SWITCH8 = 0, JTAG CONNECTOR WHEN SWITCH8 = 1
--
JTAG_TCK			<= USBC_0 WHEN SWITCH8 = '0' ELSE 'Z';
JTAG_TDI			<= USBC_1 WHEN SWITCH8 = '0' ELSE 'Z';
USBC_2			<= JTAG_TDO;
JTAG_TMS			<= USBC_3 WHEN SWITCH8 = '0' ELSE 'Z';
-- SPI Signals driven from USB Port 1 when SWITCH6 = 1, DETACHED WHEN SWITCH6 = 0
SPI_SK			<= USBC_8 WHEN SWITCH6 = '1' ELSE 'Z';
SPI_DO			<= USBC_9 WHEN SWITCH6 = '1' ELSE 'Z';
USBC_10			<= SPI_DI;
SPI_CS			<= USBC_11 WHEN SWITCH6 = '1' ELSE 'Z';
--
-- Control Power Supplies for each Array FPGA
--
--
-- SWITCH3 NOW STOPS THE CLOCK ALSO TO THE ARRAY
--
--was CLOCK_STOP 		<= SWITCH8 OR SWITCH3;
CLOCK_STOP 		<= SWITCH3;
--
-- SWITCH4 - SET LOOPBACK ON FOR UP-LINK AND DOWN-LINK 4 BITS EACH
--
LBACK: LOOPBACK_TEST		
	PORT MAP(
		CLOCK_50MHZ       => 	CLOCK_25MHZ,
      RESET_N 		      => 	RESET_N,
      IO_TEST_BUS_IN(1)	=>		LOOPIN1,
		IO_TEST_BUS_IN(2)	=>		LOOPIN2,
		IO_TEST_BUS_IN(3)	=>		LOOPIN3,
		IO_TEST_BUS_IN(4)	=>		LOOPIN4,
      IO_TEST_BUS_OUT(1)=>		LOOPOUT1,
      IO_TEST_BUS_OUT(2)=>		LOOPOUT2,
      IO_TEST_BUS_OUT(3)=>		LOOPOUT3,
      IO_TEST_BUS_OUT(4)=>		LOOPOUT4,
		LOOPBACK_PASS  	=> 	LOOPBACK_PASS
		);
--
-- ENABLE LOOPBACKS WHEN SWITCH4 = 1
--
      LOOPIN1		<= UP1 WHEN SWITCH4 = '1' ELSE '0';
		LOOPIN2		<= UP2 WHEN SWITCH4 = '1' ELSE '0';
		LOOPIN3		<= UP3 WHEN SWITCH4 = '1' ELSE '0';
		LOOPIN4		<= UP4 WHEN SWITCH4 = '1' ELSE '0';
      DOWN1 	   <= LOOPOUT1 WHEN SWITCH4 = '1' ELSE 'Z';
      DOWN2   	   <= LOOPOUT2 WHEN SWITCH4 = '1' ELSE 'Z';
      DOWN3	      <= LOOPOUT3 WHEN SWITCH4 = '1' ELSE 'Z';
      DOWN4	      <= LOOPOUT4 WHEN SWITCH4 = '1' ELSE 'Z';
		LED			<= FLASH WHEN SWITCH4 = '0' ELSE LOOPBACK_PASS;
--
-- ENABLE THE 3V3 WHEN ANY OF THE 1V2'S ARE ENABLED
--
--ARRAY_3V3_EN 	<= '0' WHEN ((SWITCH1 = '0') OR (SWITCH2 = '0') OR (SWITCH3 = '0') OR (SWITCH4 = '0')) ELSE '1';
--
-- ROUTE TX,RX FROM FTDI PORT 2 & 3 (0 IS DEDICATED JTAG FOR ARRAY, 1 IS DEDICATED SPI FOR 3S50AN)
--
-- FPGA 1
USB1_1			<= USBC_16; -- TXD (OUT)
USBC_17			<= USB1_2;  -- RXD (IN)
-- FPGA 3
USB3_1			<= USBC_24;	-- TXD (OUT)
USBC_25			<= USB3_2;	-- RXD (IN)
--
--




divide1 : PROCESS(RESET,CLK50)
BEGIN
IF (RESET = '1') THEN
   CLOCK_DIVIDE_COUNTER <= 24999; 
   TOGGLE_1KHZ          <= '0';  
   CLOCK_1KHZ           <= '0';    
   
ELSIF (CLK50'event  AND CLK50='1') THEN
   IF (CLOCK_DIVIDE_COUNTER = 0) THEN
      CLOCK_DIVIDE_COUNTER <= 24999; 
      TOGGLE_1KHZ          <= '1';  
   ELSE
      CLOCK_DIVIDE_COUNTER <= CLOCK_DIVIDE_COUNTER -1; 
      TOGGLE_1KHZ          <= '0';  
   END IF;
   
   IF (TOGGLE_1KHZ = '1') THEN
      IF (CLOCK_1KHZ = '1') THEN
         CLOCK_1KHZ <= '0';    
      ELSE
         CLOCK_1KHZ <= '1';    
      END IF;
   ELSE
      CLOCK_1KHZ <= CLOCK_1KHZ;   
   END IF;
   
   
   
END IF;
END PROCESS divide1;





INDICATOR1 : PROCESS(SWITCH5)
BEGIN
   IF (SWITCH5 ='1') THEN
      FREQUENCY_IS_100MHZ <= '1'; 
   ELSE
      FREQUENCY_IS_100MHZ <= '0'; 
   END IF;

   IF (SWITCH5 ='0') THEN
      FREQUENCY_IS_50MHZ <= '1'; 
   ELSE
      FREQUENCY_IS_50MHZ <= '0'; 
   END IF;
   
   
   
END PROCESS INDICATOR1;


CLKOP : PROCESS(CLK50)
BEGIN
IF (CLK50'event  AND CLK50='1') THEN
	USB1_5   <= CLOCK_1KHZ;
	USB2_5	<= CLOCK_1KHZ;
	USB3_5	<= CLOCK_1KHZ;
	USB4_5	<= CLOCK_1KHZ;


	USB1_6   <= RESET_N;
	USB2_6	<= RESET_N;
	USB3_6	<= RESET_N;
	USB4_6	<= RESET_N;


	USB1_7   <= FREQUENCY_IS_100MHZ;
	USB2_7	<= FREQUENCY_IS_100MHZ;
	USB3_7	<= FREQUENCY_IS_100MHZ;
	USB4_7	<= FREQUENCY_IS_100MHZ;

END IF;
END PROCESS CLKOP;




TURNON : PROCESS(RESET,CLOCK_25MHZ)
BEGIN
IF (RESET = '1') THEN
   COUNTER_100MS        <= 24999999;
   COUNTER_100MS_TICK   <= '0';
   POWER_STARTUP_N      <= "111111";

ELSIF (CLOCK_25MHZ'EVENT  AND CLOCK_25MHZ='1') THEN
   IF (POWER_STARTUP_N(5) = '1') THEN
      IF (COUNTER_100MS = 0) THEN
         COUNTER_100MS        <= 24999999;
         COUNTER_100MS_TICK   <= '1';
      ELSE
         COUNTER_100MS        <= COUNTER_100MS - 1;
         COUNTER_100MS_TICK   <= '0';
      END IF;
   ELSE
      COUNTER_100MS        <= 24999999;
      COUNTER_100MS_TICK   <= '0';
   END IF;

   
   --NO FAN = NO 12V OR OVERRIDDEN
   IF (FAN_IS_RUNNING = '0') THEN
      POWER_STARTUP_N(5 DOWNTO 0) <= "111111";
   --TURN THEM ON AT 100MS INTERVALS   
   ELSIF (COUNTER_100MS_TICK = '1') THEN
      POWER_STARTUP_N(5 DOWNTO 0) <= POWER_STARTUP_N(4 DOWNTO 0) & '0'; 
   --WAIT     
   ELSE
      POWER_STARTUP_N(5 DOWNTO 0) <= POWER_STARTUP_N(5 DOWNTO 0);
   END IF;

   
END IF;
END PROCESS TURNON;

ARRAY_3V3_EN	<= POWER_STARTUP_N(0);     -- ON = SUPPLY ON
EN_1V2_1			<= POWER_STARTUP_N(1);		-- ON = SUPPLY ON
EN_1V2_2			<= POWER_STARTUP_N(2);		-- ON = SUPPLY ON
EN_1V2_3			<= POWER_STARTUP_N(3);		-- ON = SUPPLY ON
EN_1V2_4			<= POWER_STARTUP_N(4);		-- ON = SUPPLY ON



FAN1 : PROCESS(RESET,CLOCK_25MHZ)
BEGIN
IF (RESET = '1') THEN
   TICK_COUNTER         <=  0 ;
   TICK_1SEC            <= '0';
   FAN_RPM1_SHIFT       <= (OTHERS => '0');
   FAN_RPM2_SHIFT       <= (OTHERS => '0');
   FAN_RPM3_SHIFT       <= (OTHERS => '0');
   FAN_RPM4_SHIFT       <= (OTHERS => '0');
   FAN_COUNTER1         <= (OTHERS => '0');
   FAN_COUNTER2         <= (OTHERS => '0');
   FAN_COUNTER3         <= (OTHERS => '0');
   FAN_COUNTER4         <= (OTHERS => '0');
   FAN_COUNTER1_STORED  <= (OTHERS => '0');
   FAN_COUNTER2_STORED  <= (OTHERS => '0');
   FAN_COUNTER3_STORED  <= (OTHERS => '0');
   FAN_COUNTER4_STORED  <= (OTHERS => '0');
   FAN1_IS_OK           <= '0';
   FAN2_IS_OK           <= '0';
   FAN3_IS_OK           <= '0';
   FAN4_IS_OK           <= '0';
   FAN_IS_RUNNING       <= '0';
   
ELSIF (CLOCK_25MHZ'EVENT  AND CLOCK_25MHZ='1') THEN
   IF (TICK_COUNTER = 0) THEN
      TICK_COUNTER <= 24999999;   
      TICK_1SEC    <= '1';
   ELSE
      TICK_COUNTER <= TICK_COUNTER - 1;   
      TICK_1SEC    <= '0';
   END IF;

   FAN_RPM1_SHIFT <= FAN_RPM1_SHIFT(2 downto 0) & FAN_RPM1;
   FAN_RPM2_SHIFT <= FAN_RPM2_SHIFT(2 downto 0) & FAN_RPM2;
   FAN_RPM3_SHIFT <= FAN_RPM3_SHIFT(2 downto 0) & FAN_RPM3;
   FAN_RPM4_SHIFT <= FAN_RPM4_SHIFT(2 downto 0) & FAN_RPM4;

   IF    (TICK_1SEC = '1') THEN
      FAN_COUNTER1   <= (OTHERS => '0');
   ELSIF (FAN_RPM1_SHIFT(3 DOWNTO 2) = "01") THEN
      FAN_COUNTER1 <= FAN_COUNTER1 + 1;      
   ELSE
      FAN_COUNTER1 <= FAN_COUNTER1;      
   END IF;

   IF    (TICK_1SEC = '1') THEN
      FAN_COUNTER2   <= (OTHERS => '0');
   ELSIF (FAN_RPM2_SHIFT(3 DOWNTO 2) = "01") THEN
      FAN_COUNTER2 <= FAN_COUNTER2 + 1;      
   ELSE
      FAN_COUNTER2 <= FAN_COUNTER2;      
   END IF;

   IF    (TICK_1SEC = '1') THEN
      FAN_COUNTER3   <= (OTHERS => '0');
   ELSIF (FAN_RPM3_SHIFT(3 DOWNTO 2) = "01") THEN
      FAN_COUNTER3 <= FAN_COUNTER3 + 1;      
   ELSE
      FAN_COUNTER3 <= FAN_COUNTER3;      
   END IF;

   IF    (TICK_1SEC = '1') THEN
      FAN_COUNTER4   <= (OTHERS => '0');
   ELSIF (FAN_RPM4_SHIFT(3 DOWNTO 2) = "01") THEN
      FAN_COUNTER4 <= FAN_COUNTER4 + 1;      
   ELSE
      FAN_COUNTER4 <= FAN_COUNTER4;      
   END IF;

   IF    (TICK_1SEC = '1') THEN
      FAN_COUNTER1_STORED   <= FAN_COUNTER1;
      FAN_COUNTER2_STORED   <= FAN_COUNTER2;
      FAN_COUNTER3_STORED   <= FAN_COUNTER3;
      FAN_COUNTER4_STORED   <= FAN_COUNTER4;
   ELSE
      FAN_COUNTER1_STORED   <= FAN_COUNTER1_STORED;
      FAN_COUNTER2_STORED   <= FAN_COUNTER2_STORED;
      FAN_COUNTER3_STORED   <= FAN_COUNTER3_STORED;
      FAN_COUNTER4_STORED   <= FAN_COUNTER4_STORED;
   END IF;
   
   IF (FAN_COUNTER1_STORED(15 DOWNTO 0) > X"0017") THEN
      FAN1_IS_OK <= '1';   
   ELSE
      FAN1_IS_OK <= '0';
   END IF;

   IF (FAN_COUNTER2_STORED(15 DOWNTO 0) > X"0017") THEN
      FAN2_IS_OK <= '1';   
   ELSE
      FAN2_IS_OK <= '0';
   END IF;

   IF (FAN_COUNTER3_STORED(15 DOWNTO 0) > X"0017") THEN
      FAN3_IS_OK <= '1';   
   ELSE
      FAN3_IS_OK <= '0';
   END IF;

   IF (FAN_COUNTER4_STORED(15 DOWNTO 0) > X"0017") THEN
      FAN4_IS_OK <= '1';   
   ELSE
      FAN4_IS_OK <= '0';
   END IF;
   
   IF ((FAN1_IS_OK = '1') OR (FAN2_IS_OK = '1') OR (FAN3_IS_OK = '1') OR (FAN4_IS_OK = '1') OR (SWITCH2 = '1')) THEN
      FAN_IS_RUNNING <= '1';   
   ELSE
      FAN_IS_RUNNING <= '0';   
   END IF;


END IF;
END PROCESS FAN1;


END RTL;




